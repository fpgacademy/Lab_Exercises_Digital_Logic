
... put your processor code here
