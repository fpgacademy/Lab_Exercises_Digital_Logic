-- use your processor from Part 1

