... use your processor code from Part III

