... use your Verilog file from Part IV
