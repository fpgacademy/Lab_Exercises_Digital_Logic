... use your processor code from Part III, and add support for b{cond}
